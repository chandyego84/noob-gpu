/*
`timescale 1ns/1ps
`include "common_defs.v"

module SimdController # (

)
(

);

endmodule
*/